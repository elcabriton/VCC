module fibonacci(cvb 